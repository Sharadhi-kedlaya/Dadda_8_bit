`timescale 1ns / 1ps

module Dedda_mul(a,b,op);

input  [7:0] a,b;
output [15:0] op;

wire [7:0] p0,p1,p2,p3,p4,p5,p6,p7;

// ---------------- Partial Products ----------------
partial_product pp1(a[0],b,p0[0],p0[1],p0[2],p0[3],p0[4],p0[5],p0[6],p0[7]);
partial_product pp2(a[1],b,p1[0],p1[1],p1[2],p1[3],p1[4],p1[5],p1[6],p1[7]);
partial_product pp3(a[2],b,p2[0],p2[1],p2[2],p2[3],p2[4],p2[5],p2[6],p2[7]);
partial_product pp4(a[3],b,p3[0],p3[1],p3[2],p3[3],p3[4],p3[5],p3[6],p3[7]);
partial_product pp5(a[4],b,p4[0],p4[1],p4[2],p4[3],p4[4],p4[5],p4[6],p4[7]);
partial_product pp6(a[5],b,p5[0],p5[1],p5[2],p5[3],p5[4],p5[5],p5[6],p5[7]);
partial_product pp7(a[6],b,p6[0],p6[1],p6[2],p6[3],p6[4],p6[5],p6[6],p6[7]);
partial_product pp8(a[7],b,p7[0],p7[1],p7[2],p7[3],p7[4],p7[5],p7[6],p7[7]);

// ---------------- Intermediate Wires ----------------

wire [14:1] s1, c1;   // Level 1
wire [15:1] s2, c2;   // Level 2
wire [10:1] s3, c3;   // Level 3
wire [12:1] s4, c4;   // Level 4
wire [14:1] s5, c5;   // Level 5
wire Sf, Cf;      // Final

// ---------------- Level 1 ----------------
ha h1(p0[6],p1[5],s1[1],c1[1]);
FA f1(p0[7],p1[6],p2[5],s1[2],c1[2]);
FA f2(p1[7],p2[6],p3[5],s1[3],c1[3]);
FA f3(p2[7],p3[6],p4[5],s1[4],c1[4]);

ha h2(p3[4],p4[3],s1[5],c1[5]);
ha h3(p4[4],p5[3],s1[6],c1[6]);

// ---------------- Level 2 ----------------
ha h4(p0[4],p1[3],s2[1],c2[1]);
FA f4(p0[5],p1[4],p2[3],s2[2],c2[2]);
FA f5(s1[1],p2[4],p3[3],s2[3],c2[3]);
FA f6(s1[2],c1[1],s1[5],s2[4],c2[4]);
FA f7(s1[3],c1[2],s1[6],s2[5],c2[5]);
FA f8(s1[4],c1[3],c1[6],s2[6],c2[6]);
FA f9(c1[4],p3[7],p4[6],s2[7],c2[7]);
FA f10(p4[7],p5[6],p6[5],s2[8],c2[8]);

ha h5(p3[2],p4[1],s2[9],c2[9]);
FA f11(p4[2],p5[1],p6[0],s2[10],c2[10]);
FA f12(p5[2],p6[1],p7[0],s2[11],c2[11]);
FA f13(c1[5],p6[2],p7[1],s2[12],c2[12]);
FA f14(p5[4],p6[3],p7[2],s2[13],c2[13]);
FA f15(p5[5],p6[4],p7[3],s2[14],c2[14]);

// ---------------- Level 3 ----------------
ha h6(p0[3],p1[2],s3[1],c3[1]);
FA f16(s2[1],p2[2],p3[1],s3[2],c3[2]);
FA f17(s2[2],c2[1],s2[9],s3[3],c3[3]);
FA f18(s2[3],c2[2],c2[9],s3[4],c3[4]);
FA f19(s2[4],c2[3],s2[10],s3[5],c3[5]);
FA f20(s2[5],c2[4],s2[11],s3[6],c3[6]);
FA f21(s2[6],c2[5],s2[12],s3[7],c3[7]);
FA f22(s2[7],c2[6],s2[13],s3[8],c3[8]);
FA f23(s2[8],c2[7],p7[4],s3[9],c3[9]);
FA f24(c2[8],p5[7],p6[6],s3[10],c3[10]);

// ---------------- Level 4 ----------------
ha h7(p0[2],p1[1],s4[1],c4[1]);
FA f25(s3[1],p2[1],p3[0],s4[2],c4[2]);
FA f26(s3[2],c3[1],p4[0],s4[3],c4[3]);
FA f27(s3[3],c3[2],p5[0],s4[4],c4[4]);
FA f28(s3[4],c3[3],s2[10],s4[5],c4[5]);
FA f29(s3[5],c3[4],s2[11],s4[6],c4[6]);
FA f30(s3[6],c3[5],s2[12],s4[7],c4[7]);
FA f31(s3[7],c3[6],s2[13],s4[8],c4[8]);
FA f32(s3[8],c3[7],s2[14],s4[9],c4[9]);
FA f33(s3[9],c3[8],c2[14],s4[10],c4[10]);
FA f34(s3[10],c3[9],p7[5],s4[11],c4[11]);
FA f35(c3[10],p7[6],p6[7],s4[12],c4[12]);

// ---------------- Level 5 ----------------
ha h8(p0[1],p1[0],s5[1],c5[1]);
FA f36(s4[1],p2[0],c5[1],s5[2],c5[2]);
FA f37(s4[2],c4[1],c5[2],s5[3],c5[3]);
FA f38(s4[3],c4[2],c5[3],s5[4],c5[4]);
FA f39(s4[4],c4[3],c5[4],s5[5],c5[5]);
FA f40(s4[5],c4[4],c5[5],s5[6],c5[6]);
FA f41(s4[6],c4[5],c5[6],s5[7],c5[7]);
FA f42(s4[7],c4[6],c5[7],s5[8],c5[8]);
FA f43(s4[8],c4[7],c5[8],s5[9],c5[9]);
FA f44(s4[9],c4[8],c5[9],s5[10],c5[10]);
FA f45(s4[10],c4[9],c5[10],s5[11],c5[11]);
FA f46(s4[11],c4[10],c5[11],s5[12],c5[12]);
FA f47(s4[12],c4[11],c5[12],s5[13],c5[13]);
  FA f48(p7[7],c4[12],c5[13],Sf,Cf);

// ---------------- Final Output ----------------
  assign op = {Cf,Sf,s5[13],s5[12],s5[11],s5[10],
             s5[9],s5[8],s5[7],s5[6],s5[5],s5[4],
             s5[3],s5[2],s5[1],p0[0]};

endmodule

